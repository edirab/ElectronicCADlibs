UA741 OPAMP
.OPTIONS ACCT
.OP
*ALIAS V(6)=VOUT
*ALIAS V(2)=VSUM
Q6 24 12 21 QNL
R14 13 4 1K
R2 21 4 1K
Q7 20 16 12 QNL
R3 12 4 50K
Q24 16 15 3 QPL
Q4 24 15 25 QPL
Q1 10 0 3 QNL
Q2 10 2 25 QNL
Q10 10 10 20 QPL
Q11 15 10 20 QPL
Q8 15 23 9 QNL
Q9 23 23 4 QNL
R4 9 4 5K
Q12 18 18 20 QPL
Q18 19 24 14 QNL
Q19 19 14 11 QNL
R5 11 4 100
Q13 24 31 4 QNL
R6 14 4 50K
Q14 5 18 20 QPL
Q15 5 8 19 QNL
R7 8 5 50K
R8 8 19 50K
R9 18 23 39K
C2 5 24 30P
Q20 5 26 6 QNL
Q22 20 5 26 QNL
R10 26 6 50
R11 6 17 25
Q23 4 19 17 QPL
V3 0 4 15
V2 20 0 15
R12 2 1 100K
V4 1 0 PULSE 0 5 0 0 0 25U
R13 2 6 100K
Q21 31 17 6 QPL
Q17 31 31 4 QNL
C3 6 0 15P
Q3 16 12 13 QNL
   .MODEL QNL NPN BF=80 RB=100 CCS=2PF TF=0.3NS TR=6NS CJE=3PF CJC=2PF VAF=50
   .MODEL QPL PNP BF=10 RB=20 TF=1NS TR=20NS CJE=6PF CJC=4PF VAF=50
*.PROBE
.TRAN 2.5e-007 50U 0 0
.TEMP 27
.PLOT TRAN V(6) 0.4,-5.5
.PLOT TRAN V(2) 3,-3
.PRINT TRAN V(6) V(2) 
.END
