rtlinv
*SPICE_NET
.MODEL QND NPN BF=50 RB=70 RC=40 CCS=2PF TF=0.1NS TR=10NS
+ CJE=0.9PF CJC=1.5PF PC=0.85 VA=50
Q2 4 1 0 QND
RB1 6 5 10K
RC1 3 2 1K
RC2 4 2 1K
RB2 3 1 10K
VIN 6 0 PULSE 0 5 2NS 2NS 2NS 80NS
VCC 2 0 5
Q1 3 5 0 QND
.TRAN 2e-009 200NS 0 0
.PLOT TRAN V(4) V(3) 5.5,0
.PRINT TRAN V(4) V(3) 
.AC DEC -0.5 1e+006 1e+008
.PLOT AC VM(4) VM(3) 1,-1
.PLOT AC VP(4) VP(3) 1,-1
.PRINT AC VM(4)
.PRINT AC VP(4)
.PRINT AC VM(3)
.PRINT AC VP(3)
.dc VIN 0 5 0.1
.TEMP 101
.PLOT DC V(4) V(3) 5.5,0
.PRINT DC V(4) V(3)
.END

