*jedec PLA file test
u1 stim(1,1) $g_dpwr $g_dgnd clk
+IO_STM
+0ns 0
+label=start
+50ns 1
+100ns 0
+150ns goto start -1 times

u2 stim(1,1) $g_dpwr $g_dgnd rst1
+IO_STM
+0ns 1
+60NS 0
+1000NS 0
+1500NS 0
+2000NS 0

u3 stim(1,1) $g_dpwr $g_dgnd rst2
+IO_STM
+0ns 1
+30ns 0
+1000NS 0
+2000NS 0

u3A stim(1,1) $g_dpwr $g_dgnd HI
+IO_STM
+0ns 1

X1 CLK RST1 RST2 HI HI HI HI HI HI HI
+HI HI IO1 IO2 IO5 IO6 IO9 IO10 IO8 IO7 IO4 IO3 P22V10
+  TEXT: JEDEC_FILE = "PLA1.JED"

.subckt P22V10 PIN1 PIN2 PIN3 PIN4 PIN5 PIN6 PIN7 PIN8 PIN9 PIN10 PIN11
+  PIN13 PIN14 PIN15 PIN16 PIN17 PIN18 PIN19 PIN20 PIN21 PIN22 PIN23
+  optional: PIN24=$G_DPWR PIN12=$G_DGND
+  params: MNTYMXDLY=0 IO_LEVEL=0
+  text: JEDEC_FILE="PLATEST1.JED"

U4 PLANDC(22,132) PIN24 PIN12
+  PIN1 PIN23B PIN2 PIN22B PIN3 PIN21B PIN4 PIN20B PIN5 PIN19B
+  PIN6 PIN18B PIN7 PIN17B PIN8 PIN16B PIN9 PIN15B PIN10 PIN14B
+  PIN11 PIN13
+  ROW1 ROW2 ROW3 ROW4 ROW5 ROW6 ROW7 ROW8 ROW9 ROW10
+  ROW11 ROW12 ROW13 ROW14 ROW15 ROW16 ROW17 ROW18 ROW19 ROW20
+  ROW21 ROW22 ROW23 ROW24 ROW25 ROW26 ROW27 ROW28 ROW29 ROW30
+  ROW31 ROW32 ROW33 ROW34 ROW35 ROW36 ROW37 ROW38 ROW39 ROW40
+  ROW41 ROW42 ROW43 ROW44 ROW45 ROW46 ROW47 ROW48 ROW49 ROW50
+  ROW51 ROW52 ROW53 ROW54 ROW55 ROW56 ROW57 ROW58 ROW59 ROW60
+  ROW61 ROW62 ROW63 ROW64 ROW65 ROW66 ROW67 ROW68 ROW69 ROW70
+  ROW71 ROW72 ROW73 ROW74 ROW75 ROW76 ROW77 ROW78 ROW79 ROW80
+  ROW81 ROW82 ROW83 ROW84 ROW85 ROW86 ROW87 ROW88 ROW89 ROW90
+  ROW91 ROW92 ROW93 ROW94 ROW95 ROW96 ROW97 ROW98 ROW99 ROW100
+  ROW101 ROW102 ROW103 ROW104 ROW105 ROW106 ROW107 ROW108 ROW109 ROW110
+  ROW111 ROW112 ROW113 ROW114 ROW115 ROW116 ROW117 ROW118 ROW119 ROW120
+  ROW121 ROW122 ROW123 ROW124 ROW125 ROW126 ROW127 ROW128 ROW129 ROW130
+  ROW131 ROW132
+  D0_PLD IO_LS MNTYMXDLY={MNTYMXDLY} IO_LEVEL={IO_LEVEL}
+  FILE=|JEDEC_FILE|

U5 ORA(8,2) PIN24 PIN12
+  ROW3 ROW4 ROW5 ROW6 ROW7 ROW8 ROW9 ROW10
+  ROW124 ROW125 ROW126 ROW127 ROW128 ROW129 ROW130 ROW131
+  OR1 OR10
+  D0_GATE IO_STD MNTYMXDLY={MNTYMXDLY} IO_LEVEL={IO_LEVEL}

U6 ORA(10,2) PIN24 PIN12
+  ROW12 ROW13 ROW14 ROW15 ROW16 ROW17 ROW18 ROW19 ROW20 ROW21
+  ROW113 ROW114 ROW115 ROW116 ROW117 ROW118 ROW119 ROW120 ROW121 ROW122
+  OR2 OR9
+  D0_GATE IO_STD MNTYMXDLY={MNTYMXDLY} IO_LEVEL={IO_LEVEL}

U7 ORA(12,2) PIN24 PIN12
+  ROW23 ROW24 ROW25 ROW26 ROW27 ROW28 ROW29 ROW30 ROW31 ROW32
+  ROW33 ROW34
+  ROW100 ROW101 ROW102 ROW103 ROW104 ROW105 ROW106 ROW107 ROW108 ROW109
+  ROW110 ROW111
+  OR3 OR8
+  D0_GATE IO_STD MNTYMXDLY={MNTYMXDLY} IO_LEVEL={IO_LEVEL}

U8 ORA(14,2) PIN24 PIN12
+  ROW36 ROW37 ROW38 ROW39 ROW40 ROW41 ROW42 ROW43 ROW44 ROW45
+  ROW46 ROW47 ROW48 ROW49
+  ROW85 ROW86 ROW87 ROW88 ROW89 ROW90 ROW91 ROW92 ROW93 ROW94
+  ROW95 ROW96 ROW97 ROW98
+  OR4 OR7
+  D0_GATE IO_STD MNTYMXDLY={MNTYMXDLY} IO_LEVEL={IO_LEVEL}

U9 ORA(16,2) PIN24 PIN12
+  ROW51 ROW52 ROW53 ROW54 ROW55 ROW56 ROW57 ROW58 ROW59 ROW60
+  ROW61 ROW62 ROW63 ROW64 ROW65 ROW66
+  ROW68 ROW69 ROW70 ROW71 ROW72 ROW73 ROW74 ROW75 ROW76 ROW77
+  ROW78 ROW79 ROW80 ROW81 ROW82 ROW83
+  OR5 OR6
+  D0_GATE IO_STD MNTYMXDLY={MNTYMXDLY} IO_LEVEL={IO_LEVEL}

U10A INVA(2) PIN24 PIN12
+  ROW132 ROW1 SP AR
+  D0_GATE IO_STD MNTYMXDLY={MNTYMXDLY} IO_LEVEL={IO_LEVEL}

U10 DFF(10) PIN24 PIN12
+  SP AR PIN1
+  OR1 OR2 OR3 OR4 OR5 OR6 OR7 OR8 OR9 OR10
+  P23 P22 P21 P20 P19 P18 P17 P16 P15 P14
+  PIN23B PIN22B PIN21B PIN20B PIN19B PIN18B PIN17B PIN16B PIN15B PIN14B
+  D0_EFF IO_STD MNTYMXDLY={MNTYMXDLY} IO_LEVEL={IO_LEVEL}

U11 BUF3 PIN24 PIN12
+  P23 ROW2 PIN23
+  DO_TGATE IO_STD MNTYMXDLY={MNTYMXDLY} IO_LEVEL={IO_LEVEL}

U12 BUF3 PIN24 PIN12
+  P22 ROW11 PIN22
+  DO_TGATE IO_STD MNTYMXDLY={MNTYMXDLY} IO_LEVEL={IO_LEVEL}

U13 BUF3 PIN24 PIN12
+  P21 ROW22 PIN21
+  DO_TGATE IO_STD MNTYMXDLY={MNTYMXDLY} IO_LEVEL={IO_LEVEL}

U14 BUF3 PIN24 PIN12
+  P20 ROW35 PIN20
+  DO_TGATE IO_STD MNTYMXDLY={MNTYMXDLY} IO_LEVEL={IO_LEVEL}

U15 BUF3 PIN24 PIN12
+  P19 ROW50 PIN19
+  DO_TGATE IO_STD MNTYMXDLY={MNTYMXDLY} IO_LEVEL={IO_LEVEL}

U16 BUF3 PIN24 PIN12
+  P18 ROW67 PIN18
+  DO_TGATE IO_STD MNTYMXDLY={MNTYMXDLY} IO_LEVEL={IO_LEVEL}

U17 BUF3 PIN24 PIN12
+  P17 ROW84 PIN17
+  DO_TGATE IO_STD MNTYMXDLY={MNTYMXDLY} IO_LEVEL={IO_LEVEL}

U18 BUF3 PIN24 PIN12
+  P16 ROW99 PIN16
+  DO_TGATE IO_STD MNTYMXDLY={MNTYMXDLY} IO_LEVEL={IO_LEVEL}

U19 BUF3 PIN24 PIN12
+  P15 ROW112 PIN15
+  DO_TGATE IO_STD MNTYMXDLY={MNTYMXDLY} IO_LEVEL={IO_LEVEL}

U20 BUF3 PIN24 PIN12
+  P14 ROW123 PIN14
+  DO_TGATE IO_STD MNTYMXDLY={MNTYMXDLY} IO_LEVEL={IO_LEVEL}

.ends

.MODEL DO_TGATE UTGATE ()
.MODEL D0_PLD UPLD ()

.LIB DIGIO.LIB
.PROBE
*.PRINT TRAN D(CLK) D(X1.ROW132) D(IO2) D(IO3) D(IO4) D(IO5) D(IO6) D(IO7) D(IO8) D(IO9) D(IO10) 
.TRAN 5e-008 5e-005 0 
.TEMP 27
.PLOT TRAN D(CLK) D(IO1) D(IO2) D(IO3) D(IO4) D(IO5) D(IO6) D(IO7) D(IO8) D(IO9)
+ D(IO10)
.END
