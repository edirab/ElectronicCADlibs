E:\MC7\DATA\ECLGATE.CIR Transient Analysis
* Spectrum Software Bill Steele
*
D1 13 14 D1
D2 12 15 D1
Q1 1 2 3 Q
Q2 0 4 3 Q
Q3 0 5 7 Q
Q4 3 8 9 Q
Q5 0 10 9 Q
Q6 0 13 4 Q
Q7 0 12 10 Q
Q8 0 1 Out Q
R1 11 10 2K
R2 13 0 100
R3 12 14 60
R4 2 17 50
R5 1 0 100
R6 11 Out 560
R7 11 15 720
R8 11 4 2K
R9 11 9 280
R10 11 8 820
R11 8 7 60
R12 5 6 50
V1 0 11 6V
VIN1 17 0 PULSE (-1.8 -0.8 1e-009 1e-009 0.995 0.005 2)
VIN2 6 0 PULSE (-0.8 -1.8 5e-009 1e-009 1e-009 5e-009 2e-008)
*
.MODEL Q NPN (BF=50 CJC=1.5P CJE=.9P VJC=0.85 RB=70 RC=40 VAF=50  
+ TF=100P TR=10N CJS=2P)
.MODEL D1 D (CJO=1000P VJ=800M BV=1K)
*
.OPTIONS ACCT LIST OPTS ABSTOL=1pA CHGTOL=.01pC DEFL=100u DEFW=100u DIGDRVF=2
+ DIGDRVZ=20K DIGERRDEFAULT=20 DIGERRLIMIT=10000 DIGFREQ=10GHz DIGINITSTATE=0
+ DIGIOLVL=2 DIGMNTYMX=2 DIGMNTYSCALE=0.4 DIGOVRDRV=3 DIGTYMXSCALE=1.6 GMIN=1p
+ ITL1=100 ITL2=50 ITL4=10 PIVREL=1m PIVTOL=.1p RELTOL=1m TNOM=27 TRTOL=7 VNTOL=1u
+ WIDTH=80
*
.TEMP 27
.TRAN 1.05263e-009 2e-008 0 
.PRINT TRAN V(17) V([OUT])
.PROBE
***  Parts Count
** Battery          1
** Resistor         12
** Diode            2
** NPN              8
** Pulse source     2
.END
