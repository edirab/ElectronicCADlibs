CHOKE.CKT
V1 1 0 SIN (0 100 50)
V2 0 3 SIN (0 100 50)
D1 1 2 DIO
D2 3 2 DIO
L1 4 2 5
R1 0 2 10K
R2 0 4 10K
C1 0 4 2UF
.MODEL DIO D (IS=1E-14 CJO=10PF)
.TRAN .2m 0.05 0 .2m
.TEMP 27
.PLOT TRAN V(1) V(2) V(3) V(4) -150,200
.END

